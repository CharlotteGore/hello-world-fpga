

`ifndef ASCII_ROM
`define ASCII_ROM

// module for 10-digit bitmap ROM
module ascii_rom(digit, yofs, bits);
  
  input [6:0] digit;		// char 0-128
  input [2:0] yofs;		// vertical offset (0-4)
  output reg [4:0] bits;	// output (5 bits)

  // combine {digit,yofs} into single ROM address
  wire [9:0] caseexpr = {digit,yofs};
  
  always @(*)
    case (caseexpr)/*{w:5,h:5,count:10}*/
//h20/32:  
10'b0100000000: bits = 5'b00000;
10'b0100000001: bits = 5'b00000;
10'b0100000010: bits = 5'b00000;
10'b0100000011: bits = 5'b00000;
10'b0100000100: bits = 5'b00000;
//h21/33: !
10'b0100001000: bits = 5'b00100;
10'b0100001001: bits = 5'b00100;
10'b0100001010: bits = 5'b00100;
10'b0100001011: bits = 5'b00000;
10'b0100001100: bits = 5'b00100;
//h22/34: "
10'b0100010000: bits = 5'b01010;
10'b0100010001: bits = 5'b01010;
10'b0100010010: bits = 5'b00000;
10'b0100010011: bits = 5'b00000;
10'b0100010100: bits = 5'b00000;
//h23/35: #
10'b0100011000: bits = 5'b01010;
10'b0100011001: bits = 5'b11111;
10'b0100011010: bits = 5'b01010;
10'b0100011011: bits = 5'b11111;
10'b0100011100: bits = 5'b01010;
//h24/36: $
10'b0100100000: bits = 5'b00100;
10'b0100100001: bits = 5'b00111;
10'b0100100010: bits = 5'b01100;
10'b0100100011: bits = 5'b00110;
10'b0100100100: bits = 5'b11100;
//h25/37: %
10'b0100101000: bits = 5'b11001;
10'b0100101001: bits = 5'b11010;
10'b0100101010: bits = 5'b00100;
10'b0100101011: bits = 5'b01011;
10'b0100101100: bits = 5'b10011;
//h26/38: &
10'b0100110000: bits = 5'b01000;
10'b0100110001: bits = 5'b01000;
10'b0100110010: bits = 5'b10101;
10'b0100110011: bits = 5'b10010;
10'b0100110100: bits = 5'b01101;
//h27/39: '
10'b0100111000: bits = 5'b00100;
10'b0100111001: bits = 5'b00100;
10'b0100111010: bits = 5'b00000;
10'b0100111011: bits = 5'b00000;
10'b0100111100: bits = 5'b00000;
//h28/40: (
10'b0101000000: bits = 5'b00100;
10'b0101000001: bits = 5'b01000;
10'b0101000010: bits = 5'b01000;
10'b0101000011: bits = 5'b01000;
10'b0101000100: bits = 5'b00100;
//h29/41: )
10'b0101001000: bits = 5'b00100;
10'b0101001001: bits = 5'b00010;
10'b0101001010: bits = 5'b00010;
10'b0101001011: bits = 5'b00010;
10'b0101001100: bits = 5'b00100;
//h2a/42: *
10'b0101010000: bits = 5'b10101;
10'b0101010001: bits = 5'b00100;
10'b0101010010: bits = 5'b01110;
10'b0101010011: bits = 5'b00100;
10'b0101010100: bits = 5'b10101;
//h2b/43: +
10'b0101011000: bits = 5'b00100;
10'b0101011001: bits = 5'b00100;
10'b0101011010: bits = 5'b11111;
10'b0101011011: bits = 5'b00100;
10'b0101011100: bits = 5'b00100;
//h2c/44: ,
10'b0101100000: bits = 5'b00000;
10'b0101100001: bits = 5'b00000;
10'b0101100010: bits = 5'b00000;
10'b0101100011: bits = 5'b00110;
10'b0101100100: bits = 5'b01100;
//h2d/45: -
10'b0101101000: bits = 5'b00000;
10'b0101101001: bits = 5'b00000;
10'b0101101010: bits = 5'b11111;
10'b0101101011: bits = 5'b00000;
10'b0101101100: bits = 5'b00000;
//h2e/46: .
10'b0101110000: bits = 5'b00000;
10'b0101110001: bits = 5'b00000;
10'b0101110010: bits = 5'b00000;
10'b0101110011: bits = 5'b01100;
10'b0101110100: bits = 5'b01100;
//h2f/47: /
10'b0101111000: bits = 5'b00010;
10'b0101111001: bits = 5'b00010;
10'b0101111010: bits = 5'b00100;
10'b0101111011: bits = 5'b00100;
10'b0101111100: bits = 5'b01000;
//h30/48: 0
10'b0110000000: bits = 5'b11111;
10'b0110000001: bits = 5'b10011;
10'b0110000010: bits = 5'b10101;
10'b0110000011: bits = 5'b11001;
10'b0110000100: bits = 5'b11111;
//h31/49: 1
10'b0110001000: bits = 5'b00100;
10'b0110001001: bits = 5'b01100;
10'b0110001010: bits = 5'b00100;
10'b0110001011: bits = 5'b00100;
10'b0110001100: bits = 5'b11110;
//h32/50: 2
10'b0110010000: bits = 5'b11110;
10'b0110010001: bits = 5'b00001;
10'b0110010010: bits = 5'b01111;
10'b0110010011: bits = 5'b10000;
10'b0110010100: bits = 5'b11111;
//h33/51: 3
10'b0110011000: bits = 5'b11110;
10'b0110011001: bits = 5'b00001;
10'b0110011010: bits = 5'b01111;
10'b0110011011: bits = 5'b00001;
10'b0110011100: bits = 5'b11110;
//h34/52: 4
10'b0110100000: bits = 5'b10000;
10'b0110100001: bits = 5'b10100;
10'b0110100010: bits = 5'b11111;
10'b0110100011: bits = 5'b00100;
10'b0110100100: bits = 5'b00100;
//h35/53: 5
10'b0110101000: bits = 5'b11111;
10'b0110101001: bits = 5'b10000;
10'b0110101010: bits = 5'b11110;
10'b0110101011: bits = 5'b00001;
10'b0110101100: bits = 5'b11110;
//h36/54: 6
10'b0110110000: bits = 5'b01110;
10'b0110110001: bits = 5'b10000;
10'b0110110010: bits = 5'b11110;
10'b0110110011: bits = 5'b10001;
10'b0110110100: bits = 5'b01110;
//h37/55: 7
10'b0110111000: bits = 5'b11111;
10'b0110111001: bits = 5'b00001;
10'b0110111010: bits = 5'b00010;
10'b0110111011: bits = 5'b00010;
10'b0110111100: bits = 5'b00010;
//h38/56: 8
10'b0111000000: bits = 5'b01110;
10'b0111000001: bits = 5'b10001;
10'b0111000010: bits = 5'b01110;
10'b0111000011: bits = 5'b10001;
10'b0111000100: bits = 5'b01110;
//h39/57: 9
10'b0111001000: bits = 5'b01110;
10'b0111001001: bits = 5'b10001;
10'b0111001010: bits = 5'b01111;
10'b0111001011: bits = 5'b00001;
10'b0111001100: bits = 5'b00010;
//h3a/58: :
10'b0111010000: bits = 5'b01100;
10'b0111010001: bits = 5'b01100;
10'b0111010010: bits = 5'b00000;
10'b0111010011: bits = 5'b01100;
10'b0111010100: bits = 5'b01100;
//h3b/59: ;
10'b0111011000: bits = 5'b01100;
10'b0111011001: bits = 5'b01100;
10'b0111011010: bits = 5'b00000;
10'b0111011011: bits = 5'b01100;
10'b0111011100: bits = 5'b11000;
//h3c/60: <
10'b0111100000: bits = 5'b00100;
10'b0111100001: bits = 5'b01000;
10'b0111100010: bits = 5'b10000;
10'b0111100011: bits = 5'b01000;
10'b0111100100: bits = 5'b00100;
//h3d/61: =
10'b0111101000: bits = 5'b00000;
10'b0111101001: bits = 5'b11111;
10'b0111101010: bits = 5'b00000;
10'b0111101011: bits = 5'b11111;
10'b0111101100: bits = 5'b00000;
//h3e/62: >
10'b0111110000: bits = 5'b01000;
10'b0111110001: bits = 5'b00100;
10'b0111110010: bits = 5'b00010;
10'b0111110011: bits = 5'b00100;
10'b0111110100: bits = 5'b01000;
//h3f/63: ?
10'b0111111000: bits = 5'b11110;
10'b0111111001: bits = 5'b00001;
10'b0111111010: bits = 5'b01110;
10'b0111111011: bits = 5'b00000;
10'b0111111100: bits = 5'b01100;
//h40/64: @
10'b1000000000: bits = 5'b11111;
10'b1000000001: bits = 5'b10001;
10'b1000000010: bits = 5'b10101;
10'b1000000011: bits = 5'b10111;
10'b1000000100: bits = 5'b10000;
//h41/65: A
10'b1000001000: bits = 5'b01110;
10'b1000001001: bits = 5'b10001;
10'b1000001010: bits = 5'b11111;
10'b1000001011: bits = 5'b10001;
10'b1000001100: bits = 5'b10001;
//h42/66: B
10'b1000010000: bits = 5'b11110;
10'b1000010001: bits = 5'b10001;
10'b1000010010: bits = 5'b11111;
10'b1000010011: bits = 5'b10001;
10'b1000010100: bits = 5'b11111;
//h43/67: C
10'b1000011000: bits = 5'b11111;
10'b1000011001: bits = 5'b10000;
10'b1000011010: bits = 5'b10000;
10'b1000011011: bits = 5'b10000;
10'b1000011100: bits = 5'b11111;
//h44/68: D
10'b1000100000: bits = 5'b11110;
10'b1000100001: bits = 5'b10001;
10'b1000100010: bits = 5'b10001;
10'b1000100011: bits = 5'b10001;
10'b1000100100: bits = 5'b11111;
//h45/69: E
10'b1000101000: bits = 5'b11111;
10'b1000101001: bits = 5'b10000;
10'b1000101010: bits = 5'b11110;
10'b1000101011: bits = 5'b10000;
10'b1000101100: bits = 5'b11111;
//h46/70: F
10'b1000110000: bits = 5'b11111;
10'b1000110001: bits = 5'b10000;
10'b1000110010: bits = 5'b11100;
10'b1000110011: bits = 5'b10000;
10'b1000110100: bits = 5'b10000;
//h47/71: G
10'b1000111000: bits = 5'b11111;
10'b1000111001: bits = 5'b10000;
10'b1000111010: bits = 5'b10111;
10'b1000111011: bits = 5'b10001;
10'b1000111100: bits = 5'b11111;
//h48/72: H
10'b1001000000: bits = 5'b10001;
10'b1001000001: bits = 5'b10001;
10'b1001000010: bits = 5'b11111;
10'b1001000011: bits = 5'b10001;
10'b1001000100: bits = 5'b10001;
//h49/73: I
10'b1001001000: bits = 5'b01110;
10'b1001001001: bits = 5'b00100;
10'b1001001010: bits = 5'b00100;
10'b1001001011: bits = 5'b00100;
10'b1001001100: bits = 5'b01110;
//h4a/74: J
10'b1001010000: bits = 5'b00011;
10'b1001010001: bits = 5'b00001;
10'b1001010010: bits = 5'b00001;
10'b1001010011: bits = 5'b00001;
10'b1001010100: bits = 5'b01110;
//h4b/75: K
10'b1001011000: bits = 5'b10010;
10'b1001011001: bits = 5'b10010;
10'b1001011010: bits = 5'b11100;
10'b1001011011: bits = 5'b10010;
10'b1001011100: bits = 5'b10010;
//h4c/76: L
10'b1001100000: bits = 5'b10000;
10'b1001100001: bits = 5'b10000;
10'b1001100010: bits = 5'b10000;
10'b1001100011: bits = 5'b10000;
10'b1001100100: bits = 5'b11111;
//h4d/77: M
10'b1001101000: bits = 5'b11011;
10'b1001101001: bits = 5'b10101;
10'b1001101010: bits = 5'b10101;
10'b1001101011: bits = 5'b10101;
10'b1001101100: bits = 5'b10101;
//h4e/78: N
10'b1001110000: bits = 5'b11111;
10'b1001110001: bits = 5'b10001;
10'b1001110010: bits = 5'b10001;
10'b1001110011: bits = 5'b10001;
10'b1001110100: bits = 5'b10001;
//h4f/79: O
10'b1001111000: bits = 5'b11111;
10'b1001111001: bits = 5'b10001;
10'b1001111010: bits = 5'b10001;
10'b1001111011: bits = 5'b10001;
10'b1001111100: bits = 5'b11111;
//h50/80: P
10'b1010000000: bits = 5'b11111;
10'b1010000001: bits = 5'b10001;
10'b1010000010: bits = 5'b11111;
10'b1010000011: bits = 5'b10000;
10'b1010000100: bits = 5'b10000;
//h51/81: Q
10'b1010001000: bits = 5'b11111;
10'b1010001001: bits = 5'b10001;
10'b1010001010: bits = 5'b10101;
10'b1010001011: bits = 5'b10011;
10'b1010001100: bits = 5'b11111;
//h52/82: R
10'b1010010000: bits = 5'b11111;
10'b1010010001: bits = 5'b10001;
10'b1010010010: bits = 5'b11111;
10'b1010010011: bits = 5'b10100;
10'b1010010100: bits = 5'b10010;
//h53/83: S
10'b1010011000: bits = 5'b01111;
10'b1010011001: bits = 5'b10000;
10'b1010011010: bits = 5'b0111;
10'b1010011011: bits = 5'b00001;
10'b1010011100: bits = 5'b11110;
//h54/84: T
10'b1010100000: bits = 5'b11111;
10'b1010100001: bits = 5'b00100;
10'b1010100010: bits = 5'b00100;
10'b1010100011: bits = 5'b00100;
10'b1010100100: bits = 5'b00100;
//h55/85: U
10'b1010101000: bits = 5'b10001;
10'b1010101001: bits = 5'b10001;
10'b1010101010: bits = 5'b10001;
10'b1010101011: bits = 5'b10001;
10'b1010101100: bits = 5'b11111;
//h56/86: V
10'b1010110000: bits = 5'b10001;
10'b1010110001: bits = 5'b10001;
10'b1010110010: bits = 5'b10001;
10'b1010110011: bits = 5'b01010;
10'b1010110100: bits = 5'b00100;
//h57/87: W
10'b1010111000: bits = 5'b10001;
10'b1010111001: bits = 5'b10001;
10'b1010111010: bits = 5'b10101;
10'b1010111011: bits = 5'b10101;
10'b1010111100: bits = 5'b01010;
//h58/88: X
10'b1011000000: bits = 5'b10001;
10'b1011000001: bits = 5'b01010;
10'b1011000010: bits = 5'b00100;
10'b1011000011: bits = 5'b01010;
10'b1011000100: bits = 5'b10001;
//h59/89: Y
10'b1011001000: bits = 5'b10001;
10'b1011001001: bits = 5'b01010;
10'b1011001010: bits = 5'b00100;
10'b1011001011: bits = 5'b00100;
10'b1011001100: bits = 5'b00100;
//h5a/90: Z
10'b1011010000: bits = 5'b11111;
10'b1011010001: bits = 5'b00010;
10'b1011010010: bits = 5'b00100;
10'b1011010011: bits = 5'b01000;
10'b1011010100: bits = 5'b11111;
//h5b/91: [
10'b1011011000: bits = 5'b01110;
10'b1011011001: bits = 5'b01000;
10'b1011011010: bits = 5'b01000;
10'b1011011011: bits = 5'b01000;
10'b1011011100: bits = 5'b01110;
//h5c/92: \
10'b1011100000: bits = 5'b10000;
10'b1011100001: bits = 5'b01000;
10'b1011100010: bits = 5'b00100;
10'b1011100011: bits = 5'b00010;
10'b1011100100: bits = 5'b00001;
//h5d/93: ]
10'b1011101000: bits = 5'b01110;
10'b1011101001: bits = 5'b00010;
10'b1011101010: bits = 5'b00010;
10'b1011101011: bits = 5'b00010;
10'b1011101100: bits = 5'b01110;
//h5e/94: ^
10'b1011110000: bits = 5'b00100;
10'b1011110001: bits = 5'b01010;
10'b1011110010: bits = 5'b10001;
10'b1011110011: bits = 5'b00000;
10'b1011110100: bits = 5'b00000;
//h5f/95: _
10'b1011111000: bits = 5'b00000;
10'b1011111001: bits = 5'b00000;
10'b1011111010: bits = 5'b00000;
10'b1011111011: bits = 5'b00000;
10'b1011111100: bits = 5'b11111;
//h60/96: `
10'b1100000000: bits = 5'b01100;
10'b1100000001: bits = 5'b00110;
10'b1100000010: bits = 5'b00000;
10'b1100000011: bits = 5'b00000;
10'b1100000100: bits = 5'b00000;
//h61/97: a
10'b1100001000: bits = 5'b01110;
10'b1100001001: bits = 5'b00001;
10'b1100001010: bits = 5'b01111;
10'b1100001011: bits = 5'b10001;
10'b1100001100: bits = 5'b11111;
//h62/98: b
10'b1100010000: bits = 5'b10000;
10'b1100010001: bits = 5'b11110;
10'b1100010010: bits = 5'b10001;
10'b1100010011: bits = 5'b10001;
10'b1100010100: bits = 5'b11110;
//h63/99: c
10'b1100011000: bits = 5'b00000;
10'b1100011001: bits = 5'b01110;
10'b1100011010: bits = 5'b10000;
10'b1100011011: bits = 5'b10000;
10'b1100011100: bits = 5'b01110;
//h64/100: d
10'b1100100000: bits = 5'b00001;
10'b1100100001: bits = 5'b01111;
10'b1100100010: bits = 5'b10001;
10'b1100100011: bits = 5'b10001;
10'b1100100100: bits = 5'b01111;
//h65/101: e
10'b1100101000: bits = 5'b01110;
10'b1100101001: bits = 5'b10001;
10'b1100101010: bits = 5'b11110;
10'b1100101011: bits = 5'b10000;
10'b1100101100: bits = 5'b01110;
//h66/102: f
10'b1100110000: bits = 5'b00000;
10'b1100110001: bits = 5'b00110;
10'b1100110010: bits = 5'b01000;
10'b1100110011: bits = 5'b01100;
10'b1100110100: bits = 5'b01000;
//h67/103: g
10'b1100111000: bits = 5'b11110;
10'b1100111001: bits = 5'b10010;
10'b1100111010: bits = 5'b11110;
10'b1100111011: bits = 5'b00010;
10'b1100111100: bits = 5'b11100;
//h68/104: h
10'b1101000000: bits = 5'b10000;
10'b1101000001: bits = 5'b10000;
10'b1101000010: bits = 5'b11110;
10'b1101000011: bits = 5'b10001;
10'b1101000100: bits = 5'b10001;
//h69/105: i
10'b1101001000: bits = 5'b00100;
10'b1101001001: bits = 5'b00000;
10'b1101001010: bits = 5'b00100;
10'b1101001011: bits = 5'b00100;
10'b1101001100: bits = 5'b00100;
//h6a/106: j
10'b1101010000: bits = 5'b00100;
10'b1101010001: bits = 5'b00000;
10'b1101010010: bits = 5'b00100;
10'b1101010011: bits = 5'b00100;
10'b1101010100: bits = 5'b11000;
//h6b/107: k
10'b1101011000: bits = 5'b10000;
10'b1101011001: bits = 5'b10100;
10'b1101011010: bits = 5'b11000;
10'b1101011011: bits = 5'b10100;
10'b1101011100: bits = 5'b10010;
//h6c/108: l
10'b1101100000: bits = 5'b01000;
10'b1101100001: bits = 5'b01000;
10'b1101100010: bits = 5'b01000;
10'b1101100011: bits = 5'b01000;
10'b1101100100: bits = 5'b00110;
//h6d/109: m
10'b1101101000: bits = 5'b01010;
10'b1101101001: bits = 5'b10101;
10'b1101101010: bits = 5'b10001;
10'b1101101011: bits = 5'b10001;
10'b1101101100: bits = 5'b10001;
//h6e/110: n
10'b1101110000: bits = 5'b00000;
10'b1101110001: bits = 5'b01100;
10'b1101110010: bits = 5'b10010;
10'b1101110011: bits = 5'b10010;
10'b1101110100: bits = 5'b10010;
//h6f/111: o
10'b1101111000: bits = 5'b01100;
10'b1101111001: bits = 5'b10010;
10'b1101111010: bits = 5'b10010;
10'b1101111011: bits = 5'b10010;
10'b1101111100: bits = 5'b01100;
//h70/112: p
10'b1110000000: bits = 5'b11110;
10'b1110000001: bits = 5'b10001;
10'b1110000010: bits = 5'b11110;
10'b1110000011: bits = 5'b10000;
10'b1110000100: bits = 5'b10000;
//h71/113: q
10'b1110001000: bits = 5'b01110;
10'b1110001001: bits = 5'b10010;
10'b1110001010: bits = 5'b01110;
10'b1110001011: bits = 5'b00011;
10'b1110001100: bits = 5'b00010;
//h72/114: r
10'b1110010000: bits = 5'b00110;
10'b1110010001: bits = 5'b01000;
10'b1110010010: bits = 5'b01000;
10'b1110010011: bits = 5'b01000;
10'b1110010100: bits = 5'b01000;
//h73/115: s
10'b1110011000: bits = 5'b01110;
10'b1110011001: bits = 5'b10000;
10'b1110011010: bits = 5'b01100;
10'b1110011011: bits = 5'b00010;
10'b1110011100: bits = 5'b11100;
//h74/116: t
10'b1110100000: bits = 5'b01000;
10'b1110100001: bits = 5'b11100;
10'b1110100010: bits = 5'b01000;
10'b1110100011: bits = 5'b01000;
10'b1110100100: bits = 5'b00110;
//h75/117: u
10'b1110101000: bits = 5'b10010;
10'b1110101001: bits = 5'b10010;
10'b1110101010: bits = 5'b10010;
10'b1110101011: bits = 5'b10010;
10'b1110101100: bits = 5'b01100;
//h76/118: v
10'b1110110000: bits = 5'b10001;
10'b1110110001: bits = 5'b10001;
10'b1110110010: bits = 5'b01010;
10'b1110110011: bits = 5'b01010;
10'b1110110100: bits = 5'b00100;
//h77/119: w
10'b1110111000: bits = 5'b00000;
10'b1110111001: bits = 5'b10001;
10'b1110111010: bits = 5'b10001;
10'b1110111011: bits = 5'b10101;
10'b1110111100: bits = 5'b01010;
//h78/120: x
10'b1111000000: bits = 5'b10001;
10'b1111000001: bits = 5'b01010;
10'b1111000010: bits = 5'b00100;
10'b1111000011: bits = 5'b01010;
10'b1111000100: bits = 5'b10001;
//h79/121: y
10'b1111001000: bits = 5'b01001;
10'b1111001001: bits = 5'b01001;
10'b1111001010: bits = 5'b00111;
10'b1111001011: bits = 5'b00010;
10'b1111001100: bits = 5'b01100;
//h7a/122: z
10'b1111010000: bits = 5'b00000;
10'b1111010001: bits = 5'b11110;
10'b1111010010: bits = 5'b00010;
10'b1111010011: bits = 5'b00100;
10'b1111010100: bits = 5'b11110;
//h7b/123: {
10'b1111011000: bits = 5'b00000;
10'b1111011001: bits = 5'b00000;
10'b1111011010: bits = 5'b00000;
10'b1111011011: bits = 5'b00000;
10'b1111011100: bits = 5'b00000;
//h7c/124: |
10'b1111100000: bits = 5'b00000;
10'b1111100001: bits = 5'b00000;
10'b1111100010: bits = 5'b00000;
10'b1111100011: bits = 5'b00000;
10'b1111100100: bits = 5'b00000;
//h7d/125: }
10'b1111101000: bits = 5'b00000;
10'b1111101001: bits = 5'b00000;
10'b1111101010: bits = 5'b00000;
10'b1111101011: bits = 5'b00000;
10'b1111101100: bits = 5'b00000;
//h7e/126: ~
10'b1111110000: bits = 5'b00000;
10'b1111110001: bits = 5'b00000;
10'b1111110010: bits = 5'b00000;
10'b1111110011: bits = 5'b00000;
10'b1111110100: bits = 5'b00000;

      

      default: bits = 0;
    endcase
endmodule


`endif

/*
010 0000	040	32	20	 space
010 0001	041	33	21	!
010 0010	042	34	22	"
010 0011	043	35	23	#
010 0100	044	36	24	$
010 0101	045	37	25	%
010 0110	046	38	26	&
010 0111	047	39	27	'
010 1000	050	40	28	(
010 1001	051	41	29	)
010 1010	052	42	2A	*
010 1011	053	43	2B	+
010 1100	054	44	2C	,
010 1101	055	45	2D	-
010 1110	056	46	2E	.
010 1111	057	47	2F	/
011 0000	060	48	30	0
011 0001	061	49	31	1
011 0010	062	50	32	2
011 0011	063	51	33	3
011 0100	064	52	34	4
011 0101	065	53	35	5
011 0110	066	54	36	6
011 0111	067	55	37	7
011 1000	070	56	38	8
011 1001	071	57	39	9
011 1010	072	58	3A	:
011 1011	073	59	3B	;
011 1100	074	60	3C	<
011 1101	075	61	3D	=
011 1110	076	62	3E	>
011 1111	077	63	3F	?
100 0000	100	64	40	@	`	@
100 0001	101	65	41	A
100 0010	102	66	42	B
100 0011	103	67	43	C
100 0100	104	68	44	D
100 0101	105	69	45	E
100 0110	106	70	46	F
100 0111	107	71	47	G
100 1000	110	72	48	H
100 1001	111	73	49	I
100 1010	112	74	4A	J
100 1011	113	75	4B	K
100 1100	114	76	4C	L
100 1101	115	77	4D	M
100 1110	116	78	4E	N
100 1111	117	79	4F	O
101 0000	120	80	50	P
101 0001	121	81	51	Q
101 0010	122	82	52	R
101 0011	123	83	53	S
101 0100	124	84	54	T
101 0101	125	85	55	U
101 0110	126	86	56	V
101 0111	127	87	57	W
101 1000	130	88	58	X
101 1001	131	89	59	Y
101 1010	132	90	5A	Z
101 1011	133	91	5B	[
101 1100	134	92	5C	\	~	\
101 1101	135	93	5D	]
101 1110	136	94	5E	↑	^
101 1111	137	95	5F	←	_
110 0000	140	96	60		@	`
110 0001	141	97	61		a
110 0010	142	98	62		b
110 0011	143	99	63		c
110 0100	144	100	64		d
110 0101	145	101	65		e
110 0110	146	102	66		f
110 0111	147	103	67		g
110 1000	150	104	68		h
110 1001	151	105	69		i
110 1010	152	106	6A		j
110 1011	153	107	6B		k
110 1100	154	108	6C		l
110 1101	155	109	6D		m
110 1110	156	110	6E		n
110 1111	157	111	6F		o
111 0000	160	112	70		p
111 0001	161	113	71		q
111 0010	162	114	72		r
111 0011	163	115	73		s
111 0100	164	116	74		t
111 0101	165	117	75		u
111 0110	166	118	76		v
111 0111	167	119	77		w
111 1000	170	120	78		x
111 1001	171	121	79		y
111 1010	172	122	7A		z
111 1011	173	123	7B		{
111 1100	174	124	7C	ACK	¬	|
111 1101	175	125	7D		}
111 1110	176	126	7E	ESC	|	~
*/