
`ifndef DATAROM
`define DATAROM

module datarom(clk, row, col, digit);
  input clk;
  input [4:0] row;
  input [4:0] col;
  output reg [6:0] digit;
  
  reg [6:0] bitarray[0:31][0:31]; // ROM array (32 x 32 x 7 bits)
  assign digit = bitarray[row][col];
  
  integer i, j;
  
  initial begin
    
    // clear unused array entries
    for (i = 0; i <= 32; i++)
      for (j = 0; j <= 32; j++) 
        bitarray[i][j] = 7'b0100000; 
    
    
    bitarray[0][0] = 7'h47;
bitarray[0][1] = 7'h6f;
bitarray[0][2] = 7'h72;
bitarray[0][3] = 7'h65;
bitarray[0][4] = 7'h4f;
bitarray[0][5] = 7'h53;
bitarray[0][6] = 7'h20;
bitarray[0][7] = 7'h76;
bitarray[0][8] = 7'h30;
bitarray[0][9] = 7'h2e;
bitarray[0][10] = 7'h31;
bitarray[0][11] = 7'h20;
bitarray[0][12] = 7'h32;
bitarray[0][13] = 7'h30;
bitarray[0][14] = 7'h32;
bitarray[0][15] = 7'h30;
    
    bitarray[2][0] = 7'h41;
    bitarray[2][1] = 7'h72;
    bitarray[2][2] = 7'h72;
    bitarray[2][3] = 7'h65;
    bitarray[2][4] = 7'h73;
    bitarray[2][5] = 7'h74;
    bitarray[2][6] = 7'h20;
    bitarray[2][7] = 7'h74;
    bitarray[2][8] = 7'h68;
    bitarray[2][9] = 7'h65;
    bitarray[2][10] = 7'h20;
    bitarray[2][11] = 7'h63;
    bitarray[2][12] = 7'h6f;
    bitarray[2][13] = 7'h70;
    bitarray[2][14] = 7'h73;
    bitarray[2][15] = 7'h20;
    bitarray[2][16] = 7'h74;
    bitarray[2][17] = 7'h68;
    bitarray[2][18] = 7'h61;
    bitarray[2][19] = 7'h74;
    
bitarray[3][0] = 7'h6d;
bitarray[3][1] = 7'h75;
bitarray[3][2] = 7'h72;
bitarray[3][3] = 7'h64;
bitarray[3][4] = 7'h65;
bitarray[3][5] = 7'h72;
bitarray[3][6] = 7'h65;
bitarray[3][7] = 7'h64;
bitarray[3][8] = 7'h20;
bitarray[3][9] = 7'h42;
bitarray[3][10] = 7'h72;
bitarray[3][11] = 7'h69;
bitarray[3][12] = 7'h6f;
bitarray[3][13] = 7'h6e;
bitarray[3][14] = 7'h6e;
bitarray[3][15] = 7'h61;
bitarray[3][16] = 7'h20;
bitarray[3][17] = 7'h54;
bitarray[3][18] = 7'h61;
bitarray[3][19] = 7'h79;
bitarray[3][20] = 7'h6c;
bitarray[3][21] = 7'h6f;
bitarray[3][22] = 7'h72;
  
  end
endmodule

`endif

/*
010 0000	040	32	20	 space
010 0001	041	33	21	!
010 0010	042	34	22	"
010 0011	043	35	23	#
010 0100	044	36	24	$
010 0101	045	37	25	%
010 0110	046	38	26	&
010 0111	047	39	27	'
010 1000	050	40	28	(
010 1001	051	41	29	)
010 1010	052	42	2A	*
010 1011	053	43	2B	+
010 1100	054	44	2C	,
010 1101	055	45	2D	-
010 1110	056	46	2E	.
010 1111	057	47	2F	/
011 0000	060	48	30	0
011 0001	061	49	31	1
011 0010	062	50	32	2
011 0011	063	51	33	3
011 0100	064	52	34	4
011 0101	065	53	35	5
011 0110	066	54	36	6
011 0111	067	55	37	7
011 1000	070	56	38	8
011 1001	071	57	39	9
011 1010	072	58	3A	:
011 1011	073	59	3B	;
011 1100	074	60	3C	<
011 1101	075	61	3D	=
011 1110	076	62	3E	>
011 1111	077	63	3F	?
100 0000	100	64	40	@	`	@
100 0001	101	65	41	A
100 0010	102	66	42	B
100 0011	103	67	43	C
100 0100	104	68	44	D
100 0101	105	69	45	E
100 0110	106	70	46	F
100 0111	107	71	47	G
100 1000	110	72	48	H
100 1001	111	73	49	I
100 1010	112	74	4A	J
100 1011	113	75	4B	K
100 1100	114	76	4C	L
100 1101	115	77	4D	M
100 1110	116	78	4E	N
100 1111	117	79	4F	O
101 0000	120	80	50	P
101 0001	121	81	51	Q
101 0010	122	82	52	R
101 0011	123	83	53	S
101 0100	124	84	54	T
101 0101	125	85	55	U
101 0110	126	86	56	V
101 0111	127	87	57	W
101 1000	130	88	58	X
101 1001	131	89	59	Y
101 1010	132	90	5A	Z
101 1011	133	91	5B	[
101 1100	134	92	5C	\	~	\
101 1101	135	93	5D	]
101 1110	136	94	5E	↑	^
101 1111	137	95	5F	←	_
110 0000	140	96	60		@	`
110 0001	141	97	61		a
110 0010	142	98	62		b
110 0011	143	99	63		c
110 0100	144	100	64		d
110 0101	145	101	65		e
110 0110	146	102	66		f
110 0111	147	103	67		g
110 1000	150	104	68		h
110 1001	151	105	69		i
110 1010	152	106	6A		j
110 1011	153	107	6B		k
110 1100	154	108	6C		l
110 1101	155	109	6D		m
110 1110	156	110	6E		n
110 1111	157	111	6F		o
111 0000	160	112	70		p
111 0001	161	113	71		q
111 0010	162	114	72		r
111 0011	163	115	73		s
111 0100	164	116	74		t
111 0101	165	117	75		u
111 0110	166	118	76		v
111 0111	167	119	77		w
111 1000	170	120	78		x
111 1001	171	121	79		y
111 1010	172	122	7A		z
111 1011	173	123	7B		{
111 1100	174	124	7C	ACK	¬	|
111 1101	175	125	7D		}
111 1110	176	126	7E	ESC	|	~
*/

